module percept_bank(
   input             clk,
   input             nRst,
   input             rx,
   output            tx
);

   wire   [7:0] address [255:0];

   genvar i;
   
   generate
      for (i=0; i <= 255; i=i+1)  begin: bank
         percept percept_inst (  
            .clk           (clk        ),
            .nRst          (nRst       ),
            .address       (address[i] ),
            .rx            (rx         ),
            .tx            (tx         )
         );  
      end  
   endgenerate

   // Create an address for each percept   
   assign address[0] = 0;
   assign address[1] = 1;
   assign address[2] = 2;
   assign address[3] = 3;
   assign address[4] = 4;
   assign address[5] = 5;
   assign address[6] = 6;
   assign address[7] = 7;
   assign address[8] = 8;
   assign address[9] = 9;
   assign address[10] = 10;
   assign address[11] = 11;
   assign address[12] = 12;
   assign address[13] = 13;
   assign address[14] = 14;
   assign address[15] = 15;
   assign address[16] = 16;
   assign address[17] = 17;
   assign address[18] = 18;
   assign address[19] = 19;
   assign address[20] = 20;
   assign address[21] = 21;
   assign address[22] = 22;
   assign address[23] = 23;
   assign address[24] = 24;
   assign address[25] = 25;
   assign address[26] = 26;
   assign address[27] = 27;
   assign address[28] = 28;
   assign address[29] = 29;
   assign address[30] = 30;
   assign address[31] = 31;
   assign address[32] = 32;
   assign address[33] = 33;
   assign address[34] = 34;
   assign address[35] = 35;
   assign address[36] = 36;
   assign address[37] = 37;
   assign address[38] = 38;
   assign address[39] = 39;
   assign address[40] = 40;
   assign address[41] = 41;
   assign address[42] = 42;
   assign address[43] = 43;
   assign address[44] = 44;
   assign address[45] = 45;
   assign address[46] = 46;
   assign address[47] = 47;
   assign address[48] = 48;
   assign address[49] = 49;
   assign address[50] = 50;
   assign address[51] = 51;
   assign address[52] = 52;
   assign address[53] = 53;
   assign address[54] = 54;
   assign address[55] = 55;
   assign address[56] = 56;
   assign address[57] = 57;
   assign address[58] = 58;
   assign address[59] = 59;
   assign address[60] = 60;
   assign address[61] = 61;
   assign address[62] = 62;
   assign address[63] = 63;
   assign address[64] = 64;
   assign address[65] = 65;
   assign address[66] = 66;
   assign address[67] = 67;
   assign address[68] = 68;
   assign address[69] = 69;
   assign address[70] = 70;
   assign address[71] = 71;
   assign address[72] = 72;
   assign address[73] = 73;
   assign address[74] = 74;
   assign address[75] = 75;
   assign address[76] = 76;
   assign address[77] = 77;
   assign address[78] = 78;
   assign address[79] = 79;
   assign address[80] = 80;
   assign address[81] = 81;
   assign address[82] = 82;
   assign address[83] = 83;
   assign address[84] = 84;
   assign address[85] = 85;
   assign address[86] = 86;
   assign address[87] = 87;
   assign address[88] = 88;
   assign address[89] = 89;
   assign address[90] = 90;
   assign address[91] = 91;
   assign address[92] = 92;
   assign address[93] = 93;
   assign address[94] = 94;
   assign address[95] = 95;
   assign address[96] = 96;
   assign address[97] = 97;
   assign address[98] = 98;
   assign address[99] = 99;
   assign address[100] = 100;
   assign address[101] = 101;
   assign address[102] = 102;
   assign address[103] = 103;
   assign address[104] = 104;
   assign address[105] = 105;
   assign address[106] = 106;
   assign address[107] = 107;
   assign address[108] = 108;
   assign address[109] = 109;
   assign address[110] = 110;
   assign address[111] = 111;
   assign address[112] = 112;
   assign address[113] = 113;
   assign address[114] = 114;
   assign address[115] = 115;
   assign address[116] = 116;
   assign address[117] = 117;
   assign address[118] = 118;
   assign address[119] = 119;
   assign address[120] = 120;
   assign address[121] = 121;
   assign address[122] = 122;
   assign address[123] = 123;
   assign address[124] = 124;
   assign address[125] = 125;
   assign address[126] = 126;
   assign address[127] = 127;
   assign address[128] = 128;
   assign address[129] = 129;
   assign address[130] = 130;
   assign address[131] = 131;
   assign address[132] = 132;
   assign address[133] = 133;
   assign address[134] = 134;
   assign address[135] = 135;
   assign address[136] = 136;
   assign address[137] = 137;
   assign address[138] = 138;
   assign address[139] = 139;
   assign address[140] = 140;
   assign address[141] = 141;
   assign address[142] = 142;
   assign address[143] = 143;
   assign address[144] = 144;
   assign address[145] = 145;
   assign address[146] = 146;
   assign address[147] = 147;
   assign address[148] = 148;
   assign address[149] = 149;
   assign address[150] = 150;
   assign address[151] = 151;
   assign address[152] = 152;
   assign address[153] = 153;
   assign address[154] = 154;
   assign address[155] = 155;
   assign address[156] = 156;
   assign address[157] = 157;
   assign address[158] = 158;
   assign address[159] = 159;
   assign address[160] = 160;
   assign address[161] = 161;
   assign address[162] = 162;
   assign address[163] = 163;
   assign address[164] = 164;
   assign address[165] = 165;
   assign address[166] = 166;
   assign address[167] = 167;
   assign address[168] = 168;
   assign address[169] = 169;
   assign address[170] = 170;
   assign address[171] = 171;
   assign address[172] = 172;
   assign address[173] = 173;
   assign address[174] = 174;
   assign address[175] = 175;
   assign address[176] = 176;
   assign address[177] = 177;
   assign address[178] = 178;
   assign address[179] = 179;
   assign address[180] = 180;
   assign address[181] = 181;
   assign address[182] = 182;
   assign address[183] = 183;
   assign address[184] = 184;
   assign address[185] = 185;
   assign address[186] = 186;
   assign address[187] = 187;
   assign address[188] = 188;
   assign address[189] = 189;
   assign address[190] = 190;
   assign address[191] = 191;
   assign address[192] = 192;
   assign address[193] = 193;
   assign address[194] = 194;
   assign address[195] = 195;
   assign address[196] = 196;
   assign address[197] = 197;
   assign address[198] = 198;
   assign address[199] = 199;
   assign address[200] = 200;
   assign address[201] = 201;
   assign address[202] = 202;
   assign address[203] = 203;
   assign address[204] = 204;
   assign address[205] = 205;
   assign address[206] = 206;
   assign address[207] = 207;
   assign address[208] = 208;
   assign address[209] = 209;
   assign address[210] = 210;
   assign address[211] = 211;
   assign address[212] = 212;
   assign address[213] = 213;
   assign address[214] = 214;
   assign address[215] = 215;
   assign address[216] = 216;
   assign address[217] = 217;
   assign address[218] = 218;
   assign address[219] = 219;
   assign address[220] = 220;
   assign address[221] = 221;
   assign address[222] = 222;
   assign address[223] = 223;
   assign address[224] = 224;
   assign address[225] = 225;
   assign address[226] = 226;
   assign address[227] = 227;
   assign address[228] = 228;
   assign address[229] = 229;
   assign address[230] = 230;
   assign address[231] = 231;
   assign address[232] = 232;
   assign address[233] = 233;
   assign address[234] = 234;
   assign address[235] = 235;
   assign address[236] = 236;
   assign address[237] = 237;
   assign address[238] = 238;
   assign address[239] = 239;
   assign address[240] = 240;
   assign address[241] = 241;
   assign address[242] = 242;
   assign address[243] = 243;
   assign address[244] = 244;
   assign address[245] = 245;
   assign address[246] = 246;
   assign address[247] = 247;
   assign address[248] = 248;
   assign address[249] = 249;
   assign address[250] = 250;
   assign address[251] = 251;
   assign address[252] = 252;
   assign address[253] = 253;
   assign address[254] = 254;
   assign address[255] = 255;

endmodule
